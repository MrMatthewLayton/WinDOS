Begin3
Language:    SV, 850, Swedish
Description: FreeDOS musdrivrutin
Keywords:    Mus, hjul
End
